VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_16x52_1r1w
  FOREIGN fakeram_16x52_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.203 BY 12.753 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.140 0.072 1.164 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.004 0.072 2.028 ;
    END
  END w0_wmask_in[2]
  PIN w0_wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.868 0.072 2.892 ;
    END
  END w0_wmask_in[3]
  PIN w0_wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 0.276 10.203 0.300 ;
    END
  END w0_wmask_in[4]
  PIN w0_wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 1.140 10.203 1.164 ;
    END
  END w0_wmask_in[5]
  PIN w0_wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 2.004 10.203 2.028 ;
    END
  END w0_wmask_in[6]
  PIN w0_wmask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 2.868 10.203 2.892 ;
    END
  END w0_wmask_in[7]
  PIN w0_wmask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 12.699 0.225 12.753 ;
    END
  END w0_wmask_in[8]
  PIN w0_wmask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.639 12.699 0.657 12.753 ;
    END
  END w0_wmask_in[9]
  PIN w0_wmask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.071 12.699 1.089 12.753 ;
    END
  END w0_wmask_in[10]
  PIN w0_wmask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.503 12.699 1.521 12.753 ;
    END
  END w0_wmask_in[11]
  PIN w0_wmask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.935 12.699 1.953 12.753 ;
    END
  END w0_wmask_in[12]
  PIN w0_wmask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 12.699 2.385 12.753 ;
    END
  END w0_wmask_in[13]
  PIN w0_wmask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.799 12.699 2.817 12.753 ;
    END
  END w0_wmask_in[14]
  PIN w0_wmask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.231 12.699 3.249 12.753 ;
    END
  END w0_wmask_in[15]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.732 0.072 3.756 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.596 0.072 4.620 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.460 0.072 5.484 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.324 0.072 6.348 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 3.732 10.203 3.756 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 4.596 10.203 4.620 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 5.460 10.203 5.484 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 6.324 10.203 6.348 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.783 0.000 0.801 0.054 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.359 0.000 1.377 0.054 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.935 0.000 1.953 0.054 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.511 0.000 2.529 0.054 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.087 0.000 3.105 0.054 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.663 0.000 3.681 0.054 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.239 0.000 4.257 0.054 ;
    END
  END w0_wd_in[15]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.815 0.000 4.833 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.391 0.000 5.409 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.967 0.000 5.985 0.054 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.543 0.000 6.561 0.054 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.119 0.000 7.137 0.054 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.695 0.000 7.713 0.054 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.271 0.000 8.289 0.054 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 0.000 8.865 0.054 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.663 12.699 3.681 12.753 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.095 12.699 4.113 12.753 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 12.699 4.545 12.753 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.959 12.699 4.977 12.753 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.391 12.699 5.409 12.753 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.823 12.699 5.841 12.753 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.255 12.699 6.273 12.753 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 12.699 6.705 12.753 ;
    END
  END r0_rd_out[15]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.188 0.072 7.212 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.052 0.072 8.076 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.916 0.072 8.940 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 7.188 10.203 7.212 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 8.052 10.203 8.076 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 8.916 10.203 8.940 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.780 0.072 9.804 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.644 0.072 10.668 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.508 0.072 11.532 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 9.780 10.203 9.804 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 10.644 10.203 10.668 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 11.508 10.203 11.532 ;
    END
  END r0_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.119 12.699 7.137 12.753 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.551 12.699 7.569 12.753 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.983 12.699 8.001 12.753 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.415 12.699 8.433 12.753 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 12.699 8.865 12.753 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 10.203 12.753 ;
    LAYER M2 ;
    RECT 0 0 10.203 12.753 ;
    LAYER M3 ;
    RECT 0 0 10.203 12.753 ;
    LAYER M4 ;
    RECT 0 0 10.203 12.753 ;
  END
END fakeram_16x52_1r1w

END LIBRARY
