VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_18x256_1r1w
  FOREIGN fakeram_18x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.203 BY 46.937 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.964 0.072 2.988 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.652 0.072 5.676 ;
    END
  END w0_wmask_in[2]
  PIN w0_wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.340 0.072 8.364 ;
    END
  END w0_wmask_in[3]
  PIN w0_wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.028 0.072 11.052 ;
    END
  END w0_wmask_in[4]
  PIN w0_wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 0.276 10.203 0.300 ;
    END
  END w0_wmask_in[5]
  PIN w0_wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 2.964 10.203 2.988 ;
    END
  END w0_wmask_in[6]
  PIN w0_wmask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 5.652 10.203 5.676 ;
    END
  END w0_wmask_in[7]
  PIN w0_wmask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 8.340 10.203 8.364 ;
    END
  END w0_wmask_in[8]
  PIN w0_wmask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 46.883 0.225 46.937 ;
    END
  END w0_wmask_in[9]
  PIN w0_wmask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.603 46.883 0.621 46.937 ;
    END
  END w0_wmask_in[10]
  PIN w0_wmask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.999 46.883 1.017 46.937 ;
    END
  END w0_wmask_in[11]
  PIN w0_wmask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.395 46.883 1.413 46.937 ;
    END
  END w0_wmask_in[12]
  PIN w0_wmask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.791 46.883 1.809 46.937 ;
    END
  END w0_wmask_in[13]
  PIN w0_wmask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.187 46.883 2.205 46.937 ;
    END
  END w0_wmask_in[14]
  PIN w0_wmask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.583 46.883 2.601 46.937 ;
    END
  END w0_wmask_in[15]
  PIN w0_wmask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.979 46.883 2.997 46.937 ;
    END
  END w0_wmask_in[16]
  PIN w0_wmask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.375 46.883 3.393 46.937 ;
    END
  END w0_wmask_in[17]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.716 0.072 13.740 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.404 0.072 16.428 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.092 0.072 19.116 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.780 0.072 21.804 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.468 0.072 24.492 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 11.028 10.203 11.052 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 13.716 10.203 13.740 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 16.404 10.203 16.428 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 19.092 10.203 19.116 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.747 0.000 0.765 0.054 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.287 0.000 1.305 0.054 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.827 0.000 1.845 0.054 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 0.000 2.385 0.054 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.907 0.000 2.925 0.054 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 0.000 3.465 0.054 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.987 0.000 4.005 0.054 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 0.000 4.545 0.054 ;
    END
  END w0_wd_in[17]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.067 0.000 5.085 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.607 0.000 5.625 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.147 0.000 6.165 0.054 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 0.000 6.705 0.054 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.227 0.000 7.245 0.054 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.767 0.000 7.785 0.054 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.307 0.000 8.325 0.054 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 0.000 8.865 0.054 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.387 0.000 9.405 0.054 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.771 46.883 3.789 46.937 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.167 46.883 4.185 46.937 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.563 46.883 4.581 46.937 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.959 46.883 4.977 46.937 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.355 46.883 5.373 46.937 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.751 46.883 5.769 46.937 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.147 46.883 6.165 46.937 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.543 46.883 6.561 46.937 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.939 46.883 6.957 46.937 ;
    END
  END r0_rd_out[17]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.156 0.072 27.180 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.844 0.072 29.868 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.532 0.072 32.556 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.220 0.072 35.244 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 21.780 10.203 21.804 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 24.468 10.203 24.492 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 27.156 10.203 27.180 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 29.844 10.203 29.868 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.908 0.072 37.932 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.596 0.072 40.620 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.284 0.072 43.308 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.972 0.072 45.996 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 32.532 10.203 32.556 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 35.220 10.203 35.244 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 37.908 10.203 37.932 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 40.596 10.203 40.620 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.335 46.883 7.353 46.937 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.731 46.883 7.749 46.937 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.127 46.883 8.145 46.937 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.523 46.883 8.541 46.937 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.919 46.883 8.937 46.937 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
      RECT 0.216 13.296 9.987 13.392 ;
      RECT 0.216 14.064 9.987 14.160 ;
      RECT 0.216 14.832 9.987 14.928 ;
      RECT 0.216 15.600 9.987 15.696 ;
      RECT 0.216 16.368 9.987 16.464 ;
      RECT 0.216 17.136 9.987 17.232 ;
      RECT 0.216 17.904 9.987 18.000 ;
      RECT 0.216 18.672 9.987 18.768 ;
      RECT 0.216 19.440 9.987 19.536 ;
      RECT 0.216 20.208 9.987 20.304 ;
      RECT 0.216 20.976 9.987 21.072 ;
      RECT 0.216 21.744 9.987 21.840 ;
      RECT 0.216 22.512 9.987 22.608 ;
      RECT 0.216 23.280 9.987 23.376 ;
      RECT 0.216 24.048 9.987 24.144 ;
      RECT 0.216 24.816 9.987 24.912 ;
      RECT 0.216 25.584 9.987 25.680 ;
      RECT 0.216 26.352 9.987 26.448 ;
      RECT 0.216 27.120 9.987 27.216 ;
      RECT 0.216 27.888 9.987 27.984 ;
      RECT 0.216 28.656 9.987 28.752 ;
      RECT 0.216 29.424 9.987 29.520 ;
      RECT 0.216 30.192 9.987 30.288 ;
      RECT 0.216 30.960 9.987 31.056 ;
      RECT 0.216 31.728 9.987 31.824 ;
      RECT 0.216 32.496 9.987 32.592 ;
      RECT 0.216 33.264 9.987 33.360 ;
      RECT 0.216 34.032 9.987 34.128 ;
      RECT 0.216 34.800 9.987 34.896 ;
      RECT 0.216 35.568 9.987 35.664 ;
      RECT 0.216 36.336 9.987 36.432 ;
      RECT 0.216 37.104 9.987 37.200 ;
      RECT 0.216 37.872 9.987 37.968 ;
      RECT 0.216 38.640 9.987 38.736 ;
      RECT 0.216 39.408 9.987 39.504 ;
      RECT 0.216 40.176 9.987 40.272 ;
      RECT 0.216 40.944 9.987 41.040 ;
      RECT 0.216 41.712 9.987 41.808 ;
      RECT 0.216 42.480 9.987 42.576 ;
      RECT 0.216 43.248 9.987 43.344 ;
      RECT 0.216 44.016 9.987 44.112 ;
      RECT 0.216 44.784 9.987 44.880 ;
      RECT 0.216 45.552 9.987 45.648 ;
      RECT 0.216 46.320 9.987 46.416 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
      RECT 0.216 13.296 9.987 13.392 ;
      RECT 0.216 14.064 9.987 14.160 ;
      RECT 0.216 14.832 9.987 14.928 ;
      RECT 0.216 15.600 9.987 15.696 ;
      RECT 0.216 16.368 9.987 16.464 ;
      RECT 0.216 17.136 9.987 17.232 ;
      RECT 0.216 17.904 9.987 18.000 ;
      RECT 0.216 18.672 9.987 18.768 ;
      RECT 0.216 19.440 9.987 19.536 ;
      RECT 0.216 20.208 9.987 20.304 ;
      RECT 0.216 20.976 9.987 21.072 ;
      RECT 0.216 21.744 9.987 21.840 ;
      RECT 0.216 22.512 9.987 22.608 ;
      RECT 0.216 23.280 9.987 23.376 ;
      RECT 0.216 24.048 9.987 24.144 ;
      RECT 0.216 24.816 9.987 24.912 ;
      RECT 0.216 25.584 9.987 25.680 ;
      RECT 0.216 26.352 9.987 26.448 ;
      RECT 0.216 27.120 9.987 27.216 ;
      RECT 0.216 27.888 9.987 27.984 ;
      RECT 0.216 28.656 9.987 28.752 ;
      RECT 0.216 29.424 9.987 29.520 ;
      RECT 0.216 30.192 9.987 30.288 ;
      RECT 0.216 30.960 9.987 31.056 ;
      RECT 0.216 31.728 9.987 31.824 ;
      RECT 0.216 32.496 9.987 32.592 ;
      RECT 0.216 33.264 9.987 33.360 ;
      RECT 0.216 34.032 9.987 34.128 ;
      RECT 0.216 34.800 9.987 34.896 ;
      RECT 0.216 35.568 9.987 35.664 ;
      RECT 0.216 36.336 9.987 36.432 ;
      RECT 0.216 37.104 9.987 37.200 ;
      RECT 0.216 37.872 9.987 37.968 ;
      RECT 0.216 38.640 9.987 38.736 ;
      RECT 0.216 39.408 9.987 39.504 ;
      RECT 0.216 40.176 9.987 40.272 ;
      RECT 0.216 40.944 9.987 41.040 ;
      RECT 0.216 41.712 9.987 41.808 ;
      RECT 0.216 42.480 9.987 42.576 ;
      RECT 0.216 43.248 9.987 43.344 ;
      RECT 0.216 44.016 9.987 44.112 ;
      RECT 0.216 44.784 9.987 44.880 ;
      RECT 0.216 45.552 9.987 45.648 ;
      RECT 0.216 46.320 9.987 46.416 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 10.203 46.937 ;
    LAYER M2 ;
    RECT 0 0 10.203 46.937 ;
    LAYER M3 ;
    RECT 0 0 10.203 46.937 ;
    LAYER M4 ;
    RECT 0 0 10.203 46.937 ;
  END
END fakeram_18x256_1r1w

END LIBRARY
