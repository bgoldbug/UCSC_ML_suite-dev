VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_3x64_1r1w
  FOREIGN fakeram_3x64_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.203 BY 11.602 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 0.276 10.203 0.300 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 11.548 0.225 11.602 ;
    END
  END w0_wmask_in[2]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.620 0.072 1.644 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 1.620 10.203 1.644 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[2]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.619 0.000 2.637 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.031 0.000 5.049 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.287 11.548 1.305 11.602 ;
    END
  END r0_rd_out[2]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.964 0.072 2.988 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.308 0.072 4.332 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.652 0.072 5.676 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 2.964 10.203 2.988 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 4.308 10.203 4.332 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 5.652 10.203 5.676 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.996 0.072 7.020 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.340 0.072 8.364 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.684 0.072 9.708 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 6.996 10.203 7.020 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 8.340 10.203 8.364 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 9.684 10.203 9.708 ;
    END
  END r0_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 11.548 2.385 11.602 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 11.548 3.465 11.602 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 11.548 4.545 11.602 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.607 11.548 5.625 11.602 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 11.548 6.705 11.602 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 10.203 11.602 ;
    LAYER M2 ;
    RECT 0 0 10.203 11.602 ;
    LAYER M3 ;
    RECT 0 0 10.203 11.602 ;
    LAYER M4 ;
    RECT 0 0 10.203 11.602 ;
  END
END fakeram_3x64_1r1w

END LIBRARY
