VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_20x64_2r1w
  FOREIGN fakeram_20x64_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 12.069 BY 15.505 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.044 0.072 1.068 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.812 0.072 1.836 ;
    END
  END w0_wmask_in[2]
  PIN w0_wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.580 0.072 2.604 ;
    END
  END w0_wmask_in[3]
  PIN w0_wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.348 0.072 3.372 ;
    END
  END w0_wmask_in[4]
  PIN w0_wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 0.276 12.069 0.300 ;
    END
  END w0_wmask_in[5]
  PIN w0_wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 1.044 12.069 1.068 ;
    END
  END w0_wmask_in[6]
  PIN w0_wmask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 1.812 12.069 1.836 ;
    END
  END w0_wmask_in[7]
  PIN w0_wmask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 2.580 12.069 2.604 ;
    END
  END w0_wmask_in[8]
  PIN w0_wmask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 3.348 12.069 3.372 ;
    END
  END w0_wmask_in[9]
  PIN w0_wmask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 15.451 0.225 15.505 ;
    END
  END w0_wmask_in[10]
  PIN w0_wmask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.495 15.451 0.513 15.505 ;
    END
  END w0_wmask_in[11]
  PIN w0_wmask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.783 15.451 0.801 15.505 ;
    END
  END w0_wmask_in[12]
  PIN w0_wmask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.071 15.451 1.089 15.505 ;
    END
  END w0_wmask_in[13]
  PIN w0_wmask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.359 15.451 1.377 15.505 ;
    END
  END w0_wmask_in[14]
  PIN w0_wmask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.647 15.451 1.665 15.505 ;
    END
  END w0_wmask_in[15]
  PIN w0_wmask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.935 15.451 1.953 15.505 ;
    END
  END w0_wmask_in[16]
  PIN w0_wmask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.223 15.451 2.241 15.505 ;
    END
  END w0_wmask_in[17]
  PIN w0_wmask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.511 15.451 2.529 15.505 ;
    END
  END w0_wmask_in[18]
  PIN w0_wmask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.799 15.451 2.817 15.505 ;
    END
  END w0_wmask_in[19]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.116 0.072 4.140 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.884 0.072 4.908 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.652 0.072 5.676 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.420 0.072 6.444 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.188 0.072 7.212 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 4.116 12.069 4.140 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 4.884 12.069 4.908 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 5.652 12.069 5.676 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 6.420 12.069 6.444 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 7.188 12.069 7.212 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.567 0.000 0.585 0.054 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.927 0.000 0.945 0.054 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.287 0.000 1.305 0.054 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.647 0.000 1.665 0.054 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.007 0.000 2.025 0.054 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 0.000 2.385 0.054 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.727 0.000 2.745 0.054 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.087 0.000 3.105 0.054 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 0.000 3.465 0.054 ;
    END
  END w0_wd_in[19]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.807 0.000 3.825 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.167 0.000 4.185 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 0.000 4.545 0.054 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.887 0.000 4.905 0.054 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.247 0.000 5.265 0.054 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.607 0.000 5.625 0.054 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.967 0.000 5.985 0.054 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.327 0.000 6.345 0.054 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 0.000 6.705 0.054 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.047 0.000 7.065 0.054 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.087 15.451 3.105 15.505 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.375 15.451 3.393 15.505 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.663 15.451 3.681 15.505 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.951 15.451 3.969 15.505 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.239 15.451 4.257 15.505 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 15.451 4.545 15.505 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.815 15.451 4.833 15.505 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.103 15.451 5.121 15.505 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.391 15.451 5.409 15.505 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.679 15.451 5.697 15.505 ;
    END
  END r0_rd_out[19]
  PIN r1_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.407 0.000 7.425 0.054 ;
    END
  END r1_rd_out[0]
  PIN r1_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.767 0.000 7.785 0.054 ;
    END
  END r1_rd_out[1]
  PIN r1_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.127 0.000 8.145 0.054 ;
    END
  END r1_rd_out[2]
  PIN r1_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.487 0.000 8.505 0.054 ;
    END
  END r1_rd_out[3]
  PIN r1_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 0.000 8.865 0.054 ;
    END
  END r1_rd_out[4]
  PIN r1_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.207 0.000 9.225 0.054 ;
    END
  END r1_rd_out[5]
  PIN r1_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.567 0.000 9.585 0.054 ;
    END
  END r1_rd_out[6]
  PIN r1_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.927 0.000 9.945 0.054 ;
    END
  END r1_rd_out[7]
  PIN r1_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.287 0.000 10.305 0.054 ;
    END
  END r1_rd_out[8]
  PIN r1_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.647 0.000 10.665 0.054 ;
    END
  END r1_rd_out[9]
  PIN r1_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.967 15.451 5.985 15.505 ;
    END
  END r1_rd_out[10]
  PIN r1_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.255 15.451 6.273 15.505 ;
    END
  END r1_rd_out[11]
  PIN r1_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.543 15.451 6.561 15.505 ;
    END
  END r1_rd_out[12]
  PIN r1_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.831 15.451 6.849 15.505 ;
    END
  END r1_rd_out[13]
  PIN r1_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.119 15.451 7.137 15.505 ;
    END
  END r1_rd_out[14]
  PIN r1_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.407 15.451 7.425 15.505 ;
    END
  END r1_rd_out[15]
  PIN r1_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.695 15.451 7.713 15.505 ;
    END
  END r1_rd_out[16]
  PIN r1_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.983 15.451 8.001 15.505 ;
    END
  END r1_rd_out[17]
  PIN r1_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.271 15.451 8.289 15.505 ;
    END
  END r1_rd_out[18]
  PIN r1_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.559 15.451 8.577 15.505 ;
    END
  END r1_rd_out[19]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.956 0.072 7.980 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.724 0.072 8.748 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.492 0.072 9.516 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 7.956 12.069 7.980 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 8.724 12.069 8.748 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 9.492 12.069 9.516 ;
    END
  END w0_addr_in[5]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.260 0.072 10.284 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.028 0.072 11.052 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.796 0.072 11.820 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 10.260 12.069 10.284 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 11.028 12.069 11.052 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 11.796 12.069 11.820 ;
    END
  END r0_addr_in[5]
  PIN r1_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.564 0.072 12.588 ;
    END
  END r1_addr_in[0]
  PIN r1_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.332 0.072 13.356 ;
    END
  END r1_addr_in[1]
  PIN r1_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.100 0.072 14.124 ;
    END
  END r1_addr_in[2]
  PIN r1_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 12.564 12.069 12.588 ;
    END
  END r1_addr_in[3]
  PIN r1_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 13.332 12.069 13.356 ;
    END
  END r1_addr_in[4]
  PIN r1_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 14.100 12.069 14.124 ;
    END
  END r1_addr_in[5]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 15.451 8.865 15.505 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.135 15.451 9.153 15.505 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.423 15.451 9.441 15.505 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.711 15.451 9.729 15.505 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.999 15.451 10.017 15.505 ;
    END
  END r0_clk
  PIN r1_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.287 15.451 10.305 15.505 ;
    END
  END r1_ce_in
  PIN r1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.575 15.451 10.593 15.505 ;
    END
  END r1_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 11.853 0.336 ;
      RECT 0.216 1.008 11.853 1.104 ;
      RECT 0.216 1.776 11.853 1.872 ;
      RECT 0.216 2.544 11.853 2.640 ;
      RECT 0.216 3.312 11.853 3.408 ;
      RECT 0.216 4.080 11.853 4.176 ;
      RECT 0.216 4.848 11.853 4.944 ;
      RECT 0.216 5.616 11.853 5.712 ;
      RECT 0.216 6.384 11.853 6.480 ;
      RECT 0.216 7.152 11.853 7.248 ;
      RECT 0.216 7.920 11.853 8.016 ;
      RECT 0.216 8.688 11.853 8.784 ;
      RECT 0.216 9.456 11.853 9.552 ;
      RECT 0.216 10.224 11.853 10.320 ;
      RECT 0.216 10.992 11.853 11.088 ;
      RECT 0.216 11.760 11.853 11.856 ;
      RECT 0.216 12.528 11.853 12.624 ;
      RECT 0.216 13.296 11.853 13.392 ;
      RECT 0.216 14.064 11.853 14.160 ;
      RECT 0.216 14.832 11.853 14.928 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 11.853 0.336 ;
      RECT 0.216 1.008 11.853 1.104 ;
      RECT 0.216 1.776 11.853 1.872 ;
      RECT 0.216 2.544 11.853 2.640 ;
      RECT 0.216 3.312 11.853 3.408 ;
      RECT 0.216 4.080 11.853 4.176 ;
      RECT 0.216 4.848 11.853 4.944 ;
      RECT 0.216 5.616 11.853 5.712 ;
      RECT 0.216 6.384 11.853 6.480 ;
      RECT 0.216 7.152 11.853 7.248 ;
      RECT 0.216 7.920 11.853 8.016 ;
      RECT 0.216 8.688 11.853 8.784 ;
      RECT 0.216 9.456 11.853 9.552 ;
      RECT 0.216 10.224 11.853 10.320 ;
      RECT 0.216 10.992 11.853 11.088 ;
      RECT 0.216 11.760 11.853 11.856 ;
      RECT 0.216 12.528 11.853 12.624 ;
      RECT 0.216 13.296 11.853 13.392 ;
      RECT 0.216 14.064 11.853 14.160 ;
      RECT 0.216 14.832 11.853 14.928 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 12.069 15.505 ;
    LAYER M2 ;
    RECT 0 0 12.069 15.505 ;
    LAYER M3 ;
    RECT 0 0 12.069 15.505 ;
    LAYER M4 ;
    RECT 0 0 12.069 15.505 ;
  END
END fakeram_20x64_2r1w

END LIBRARY
