VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_32x128_2r1w
  FOREIGN fakeram_32x128_2r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 12.069 BY 30.171 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.332 0.072 1.356 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.388 0.072 2.412 ;
    END
  END w0_wmask_in[2]
  PIN w0_wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.444 0.072 3.468 ;
    END
  END w0_wmask_in[3]
  PIN w0_wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.500 0.072 4.524 ;
    END
  END w0_wmask_in[4]
  PIN w0_wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.556 0.072 5.580 ;
    END
  END w0_wmask_in[5]
  PIN w0_wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.612 0.072 6.636 ;
    END
  END w0_wmask_in[6]
  PIN w0_wmask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.668 0.072 7.692 ;
    END
  END w0_wmask_in[7]
  PIN w0_wmask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 0.276 12.069 0.300 ;
    END
  END w0_wmask_in[8]
  PIN w0_wmask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 1.332 12.069 1.356 ;
    END
  END w0_wmask_in[9]
  PIN w0_wmask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 2.388 12.069 2.412 ;
    END
  END w0_wmask_in[10]
  PIN w0_wmask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 3.444 12.069 3.468 ;
    END
  END w0_wmask_in[11]
  PIN w0_wmask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 4.500 12.069 4.524 ;
    END
  END w0_wmask_in[12]
  PIN w0_wmask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 5.556 12.069 5.580 ;
    END
  END w0_wmask_in[13]
  PIN w0_wmask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 6.612 12.069 6.636 ;
    END
  END w0_wmask_in[14]
  PIN w0_wmask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 7.668 12.069 7.692 ;
    END
  END w0_wmask_in[15]
  PIN w0_wmask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 30.117 0.225 30.171 ;
    END
  END w0_wmask_in[16]
  PIN w0_wmask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.387 30.117 0.405 30.171 ;
    END
  END w0_wmask_in[17]
  PIN w0_wmask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.567 30.117 0.585 30.171 ;
    END
  END w0_wmask_in[18]
  PIN w0_wmask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.747 30.117 0.765 30.171 ;
    END
  END w0_wmask_in[19]
  PIN w0_wmask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.927 30.117 0.945 30.171 ;
    END
  END w0_wmask_in[20]
  PIN w0_wmask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.107 30.117 1.125 30.171 ;
    END
  END w0_wmask_in[21]
  PIN w0_wmask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.287 30.117 1.305 30.171 ;
    END
  END w0_wmask_in[22]
  PIN w0_wmask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.467 30.117 1.485 30.171 ;
    END
  END w0_wmask_in[23]
  PIN w0_wmask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.647 30.117 1.665 30.171 ;
    END
  END w0_wmask_in[24]
  PIN w0_wmask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.827 30.117 1.845 30.171 ;
    END
  END w0_wmask_in[25]
  PIN w0_wmask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.007 30.117 2.025 30.171 ;
    END
  END w0_wmask_in[26]
  PIN w0_wmask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.187 30.117 2.205 30.171 ;
    END
  END w0_wmask_in[27]
  PIN w0_wmask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 30.117 2.385 30.171 ;
    END
  END w0_wmask_in[28]
  PIN w0_wmask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.547 30.117 2.565 30.171 ;
    END
  END w0_wmask_in[29]
  PIN w0_wmask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.727 30.117 2.745 30.171 ;
    END
  END w0_wmask_in[30]
  PIN w0_wmask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.907 30.117 2.925 30.171 ;
    END
  END w0_wmask_in[31]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.724 0.072 8.748 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.780 0.072 9.804 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.836 0.072 10.860 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.892 0.072 11.916 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.948 0.072 12.972 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.004 0.072 14.028 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.060 0.072 15.084 ;
    END
  END w0_wd_in[6]
  PIN w0_wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.116 0.072 16.140 ;
    END
  END w0_wd_in[7]
  PIN w0_wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 8.724 12.069 8.748 ;
    END
  END w0_wd_in[8]
  PIN w0_wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 9.780 12.069 9.804 ;
    END
  END w0_wd_in[9]
  PIN w0_wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 10.836 12.069 10.860 ;
    END
  END w0_wd_in[10]
  PIN w0_wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 11.892 12.069 11.916 ;
    END
  END w0_wd_in[11]
  PIN w0_wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 12.948 12.069 12.972 ;
    END
  END w0_wd_in[12]
  PIN w0_wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 14.004 12.069 14.028 ;
    END
  END w0_wd_in[13]
  PIN w0_wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 15.060 12.069 15.084 ;
    END
  END w0_wd_in[14]
  PIN w0_wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 16.116 12.069 16.140 ;
    END
  END w0_wd_in[15]
  PIN w0_wd_in[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[16]
  PIN w0_wd_in[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.423 0.000 0.441 0.054 ;
    END
  END w0_wd_in[17]
  PIN w0_wd_in[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.639 0.000 0.657 0.054 ;
    END
  END w0_wd_in[18]
  PIN w0_wd_in[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.855 0.000 0.873 0.054 ;
    END
  END w0_wd_in[19]
  PIN w0_wd_in[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.071 0.000 1.089 0.054 ;
    END
  END w0_wd_in[20]
  PIN w0_wd_in[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.287 0.000 1.305 0.054 ;
    END
  END w0_wd_in[21]
  PIN w0_wd_in[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.503 0.000 1.521 0.054 ;
    END
  END w0_wd_in[22]
  PIN w0_wd_in[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.719 0.000 1.737 0.054 ;
    END
  END w0_wd_in[23]
  PIN w0_wd_in[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.935 0.000 1.953 0.054 ;
    END
  END w0_wd_in[24]
  PIN w0_wd_in[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.151 0.000 2.169 0.054 ;
    END
  END w0_wd_in[25]
  PIN w0_wd_in[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 0.000 2.385 0.054 ;
    END
  END w0_wd_in[26]
  PIN w0_wd_in[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.583 0.000 2.601 0.054 ;
    END
  END w0_wd_in[27]
  PIN w0_wd_in[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.799 0.000 2.817 0.054 ;
    END
  END w0_wd_in[28]
  PIN w0_wd_in[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.015 0.000 3.033 0.054 ;
    END
  END w0_wd_in[29]
  PIN w0_wd_in[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.231 0.000 3.249 0.054 ;
    END
  END w0_wd_in[30]
  PIN w0_wd_in[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 0.000 3.465 0.054 ;
    END
  END w0_wd_in[31]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.663 0.000 3.681 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.879 0.000 3.897 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.095 0.000 4.113 0.054 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.311 0.000 4.329 0.054 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 0.000 4.545 0.054 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.743 0.000 4.761 0.054 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.959 0.000 4.977 0.054 ;
    END
  END r0_rd_out[6]
  PIN r0_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.175 0.000 5.193 0.054 ;
    END
  END r0_rd_out[7]
  PIN r0_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.391 0.000 5.409 0.054 ;
    END
  END r0_rd_out[8]
  PIN r0_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.607 0.000 5.625 0.054 ;
    END
  END r0_rd_out[9]
  PIN r0_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.823 0.000 5.841 0.054 ;
    END
  END r0_rd_out[10]
  PIN r0_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.039 0.000 6.057 0.054 ;
    END
  END r0_rd_out[11]
  PIN r0_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.255 0.000 6.273 0.054 ;
    END
  END r0_rd_out[12]
  PIN r0_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.471 0.000 6.489 0.054 ;
    END
  END r0_rd_out[13]
  PIN r0_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 0.000 6.705 0.054 ;
    END
  END r0_rd_out[14]
  PIN r0_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.903 0.000 6.921 0.054 ;
    END
  END r0_rd_out[15]
  PIN r0_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.087 30.117 3.105 30.171 ;
    END
  END r0_rd_out[16]
  PIN r0_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.267 30.117 3.285 30.171 ;
    END
  END r0_rd_out[17]
  PIN r0_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.447 30.117 3.465 30.171 ;
    END
  END r0_rd_out[18]
  PIN r0_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.627 30.117 3.645 30.171 ;
    END
  END r0_rd_out[19]
  PIN r0_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.807 30.117 3.825 30.171 ;
    END
  END r0_rd_out[20]
  PIN r0_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.987 30.117 4.005 30.171 ;
    END
  END r0_rd_out[21]
  PIN r0_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.167 30.117 4.185 30.171 ;
    END
  END r0_rd_out[22]
  PIN r0_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.347 30.117 4.365 30.171 ;
    END
  END r0_rd_out[23]
  PIN r0_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 30.117 4.545 30.171 ;
    END
  END r0_rd_out[24]
  PIN r0_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.707 30.117 4.725 30.171 ;
    END
  END r0_rd_out[25]
  PIN r0_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.887 30.117 4.905 30.171 ;
    END
  END r0_rd_out[26]
  PIN r0_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.067 30.117 5.085 30.171 ;
    END
  END r0_rd_out[27]
  PIN r0_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.247 30.117 5.265 30.171 ;
    END
  END r0_rd_out[28]
  PIN r0_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.427 30.117 5.445 30.171 ;
    END
  END r0_rd_out[29]
  PIN r0_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.607 30.117 5.625 30.171 ;
    END
  END r0_rd_out[30]
  PIN r0_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.787 30.117 5.805 30.171 ;
    END
  END r0_rd_out[31]
  PIN r1_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.119 0.000 7.137 0.054 ;
    END
  END r1_rd_out[0]
  PIN r1_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.335 0.000 7.353 0.054 ;
    END
  END r1_rd_out[1]
  PIN r1_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.551 0.000 7.569 0.054 ;
    END
  END r1_rd_out[2]
  PIN r1_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.767 0.000 7.785 0.054 ;
    END
  END r1_rd_out[3]
  PIN r1_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.983 0.000 8.001 0.054 ;
    END
  END r1_rd_out[4]
  PIN r1_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.199 0.000 8.217 0.054 ;
    END
  END r1_rd_out[5]
  PIN r1_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.415 0.000 8.433 0.054 ;
    END
  END r1_rd_out[6]
  PIN r1_rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.631 0.000 8.649 0.054 ;
    END
  END r1_rd_out[7]
  PIN r1_rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 0.000 8.865 0.054 ;
    END
  END r1_rd_out[8]
  PIN r1_rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.063 0.000 9.081 0.054 ;
    END
  END r1_rd_out[9]
  PIN r1_rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.279 0.000 9.297 0.054 ;
    END
  END r1_rd_out[10]
  PIN r1_rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.495 0.000 9.513 0.054 ;
    END
  END r1_rd_out[11]
  PIN r1_rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.711 0.000 9.729 0.054 ;
    END
  END r1_rd_out[12]
  PIN r1_rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.927 0.000 9.945 0.054 ;
    END
  END r1_rd_out[13]
  PIN r1_rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.143 0.000 10.161 0.054 ;
    END
  END r1_rd_out[14]
  PIN r1_rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.359 0.000 10.377 0.054 ;
    END
  END r1_rd_out[15]
  PIN r1_rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.967 30.117 5.985 30.171 ;
    END
  END r1_rd_out[16]
  PIN r1_rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.147 30.117 6.165 30.171 ;
    END
  END r1_rd_out[17]
  PIN r1_rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.327 30.117 6.345 30.171 ;
    END
  END r1_rd_out[18]
  PIN r1_rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.507 30.117 6.525 30.171 ;
    END
  END r1_rd_out[19]
  PIN r1_rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 30.117 6.705 30.171 ;
    END
  END r1_rd_out[20]
  PIN r1_rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.867 30.117 6.885 30.171 ;
    END
  END r1_rd_out[21]
  PIN r1_rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.047 30.117 7.065 30.171 ;
    END
  END r1_rd_out[22]
  PIN r1_rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.227 30.117 7.245 30.171 ;
    END
  END r1_rd_out[23]
  PIN r1_rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.407 30.117 7.425 30.171 ;
    END
  END r1_rd_out[24]
  PIN r1_rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.587 30.117 7.605 30.171 ;
    END
  END r1_rd_out[25]
  PIN r1_rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.767 30.117 7.785 30.171 ;
    END
  END r1_rd_out[26]
  PIN r1_rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.947 30.117 7.965 30.171 ;
    END
  END r1_rd_out[27]
  PIN r1_rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.127 30.117 8.145 30.171 ;
    END
  END r1_rd_out[28]
  PIN r1_rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.307 30.117 8.325 30.171 ;
    END
  END r1_rd_out[29]
  PIN r1_rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.487 30.117 8.505 30.171 ;
    END
  END r1_rd_out[30]
  PIN r1_rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.667 30.117 8.685 30.171 ;
    END
  END r1_rd_out[31]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.172 0.072 17.196 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.228 0.072 18.252 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.284 0.072 19.308 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.340 0.072 20.364 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 17.172 12.069 17.196 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 18.228 12.069 18.252 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 19.284 12.069 19.308 ;
    END
  END w0_addr_in[6]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.396 0.072 21.420 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.452 0.072 22.476 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.508 0.072 23.532 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.564 0.072 24.588 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 20.340 12.069 20.364 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 21.396 12.069 21.420 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 22.452 12.069 22.476 ;
    END
  END r0_addr_in[6]
  PIN r1_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.620 0.072 25.644 ;
    END
  END r1_addr_in[0]
  PIN r1_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.676 0.072 26.700 ;
    END
  END r1_addr_in[1]
  PIN r1_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.732 0.072 27.756 ;
    END
  END r1_addr_in[2]
  PIN r1_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.788 0.072 28.812 ;
    END
  END r1_addr_in[3]
  PIN r1_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 23.508 12.069 23.532 ;
    END
  END r1_addr_in[4]
  PIN r1_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 24.564 12.069 24.588 ;
    END
  END r1_addr_in[5]
  PIN r1_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 11.997 25.620 12.069 25.644 ;
    END
  END r1_addr_in[6]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 8.847 30.117 8.865 30.171 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.027 30.117 9.045 30.171 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.207 30.117 9.225 30.171 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.387 30.117 9.405 30.171 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.567 30.117 9.585 30.171 ;
    END
  END r0_clk
  PIN r1_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.747 30.117 9.765 30.171 ;
    END
  END r1_ce_in
  PIN r1_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 9.927 30.117 9.945 30.171 ;
    END
  END r1_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 11.853 0.336 ;
      RECT 0.216 1.008 11.853 1.104 ;
      RECT 0.216 1.776 11.853 1.872 ;
      RECT 0.216 2.544 11.853 2.640 ;
      RECT 0.216 3.312 11.853 3.408 ;
      RECT 0.216 4.080 11.853 4.176 ;
      RECT 0.216 4.848 11.853 4.944 ;
      RECT 0.216 5.616 11.853 5.712 ;
      RECT 0.216 6.384 11.853 6.480 ;
      RECT 0.216 7.152 11.853 7.248 ;
      RECT 0.216 7.920 11.853 8.016 ;
      RECT 0.216 8.688 11.853 8.784 ;
      RECT 0.216 9.456 11.853 9.552 ;
      RECT 0.216 10.224 11.853 10.320 ;
      RECT 0.216 10.992 11.853 11.088 ;
      RECT 0.216 11.760 11.853 11.856 ;
      RECT 0.216 12.528 11.853 12.624 ;
      RECT 0.216 13.296 11.853 13.392 ;
      RECT 0.216 14.064 11.853 14.160 ;
      RECT 0.216 14.832 11.853 14.928 ;
      RECT 0.216 15.600 11.853 15.696 ;
      RECT 0.216 16.368 11.853 16.464 ;
      RECT 0.216 17.136 11.853 17.232 ;
      RECT 0.216 17.904 11.853 18.000 ;
      RECT 0.216 18.672 11.853 18.768 ;
      RECT 0.216 19.440 11.853 19.536 ;
      RECT 0.216 20.208 11.853 20.304 ;
      RECT 0.216 20.976 11.853 21.072 ;
      RECT 0.216 21.744 11.853 21.840 ;
      RECT 0.216 22.512 11.853 22.608 ;
      RECT 0.216 23.280 11.853 23.376 ;
      RECT 0.216 24.048 11.853 24.144 ;
      RECT 0.216 24.816 11.853 24.912 ;
      RECT 0.216 25.584 11.853 25.680 ;
      RECT 0.216 26.352 11.853 26.448 ;
      RECT 0.216 27.120 11.853 27.216 ;
      RECT 0.216 27.888 11.853 27.984 ;
      RECT 0.216 28.656 11.853 28.752 ;
      RECT 0.216 29.424 11.853 29.520 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 11.853 0.336 ;
      RECT 0.216 1.008 11.853 1.104 ;
      RECT 0.216 1.776 11.853 1.872 ;
      RECT 0.216 2.544 11.853 2.640 ;
      RECT 0.216 3.312 11.853 3.408 ;
      RECT 0.216 4.080 11.853 4.176 ;
      RECT 0.216 4.848 11.853 4.944 ;
      RECT 0.216 5.616 11.853 5.712 ;
      RECT 0.216 6.384 11.853 6.480 ;
      RECT 0.216 7.152 11.853 7.248 ;
      RECT 0.216 7.920 11.853 8.016 ;
      RECT 0.216 8.688 11.853 8.784 ;
      RECT 0.216 9.456 11.853 9.552 ;
      RECT 0.216 10.224 11.853 10.320 ;
      RECT 0.216 10.992 11.853 11.088 ;
      RECT 0.216 11.760 11.853 11.856 ;
      RECT 0.216 12.528 11.853 12.624 ;
      RECT 0.216 13.296 11.853 13.392 ;
      RECT 0.216 14.064 11.853 14.160 ;
      RECT 0.216 14.832 11.853 14.928 ;
      RECT 0.216 15.600 11.853 15.696 ;
      RECT 0.216 16.368 11.853 16.464 ;
      RECT 0.216 17.136 11.853 17.232 ;
      RECT 0.216 17.904 11.853 18.000 ;
      RECT 0.216 18.672 11.853 18.768 ;
      RECT 0.216 19.440 11.853 19.536 ;
      RECT 0.216 20.208 11.853 20.304 ;
      RECT 0.216 20.976 11.853 21.072 ;
      RECT 0.216 21.744 11.853 21.840 ;
      RECT 0.216 22.512 11.853 22.608 ;
      RECT 0.216 23.280 11.853 23.376 ;
      RECT 0.216 24.048 11.853 24.144 ;
      RECT 0.216 24.816 11.853 24.912 ;
      RECT 0.216 25.584 11.853 25.680 ;
      RECT 0.216 26.352 11.853 26.448 ;
      RECT 0.216 27.120 11.853 27.216 ;
      RECT 0.216 27.888 11.853 27.984 ;
      RECT 0.216 28.656 11.853 28.752 ;
      RECT 0.216 29.424 11.853 29.520 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 12.069 30.171 ;
    LAYER M2 ;
    RECT 0 0 12.069 30.171 ;
    LAYER M3 ;
    RECT 0 0 12.069 30.171 ;
    LAYER M4 ;
    RECT 0 0 12.069 30.171 ;
  END
END fakeram_32x128_2r1w

END LIBRARY
