VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_7x256_1r1w
  FOREIGN fakeram_7x256_1r1w 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.203 BY 45.963 ;
  CLASS BLOCK ;
  PIN w0_wmask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.276 0.072 0.300 ;
    END
  END w0_wmask_in[0]
  PIN w0_wmask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.020 0.072 4.044 ;
    END
  END w0_wmask_in[1]
  PIN w0_wmask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 0.276 10.203 0.300 ;
    END
  END w0_wmask_in[2]
  PIN w0_wmask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 4.020 10.203 4.044 ;
    END
  END w0_wmask_in[3]
  PIN w0_wmask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 45.909 0.225 45.963 ;
    END
  END w0_wmask_in[4]
  PIN w0_wmask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.927 45.909 0.945 45.963 ;
    END
  END w0_wmask_in[5]
  PIN w0_wmask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.647 45.909 1.665 45.963 ;
    END
  END w0_wmask_in[6]
  PIN w0_wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.764 0.072 7.788 ;
    END
  END w0_wd_in[0]
  PIN w0_wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.508 0.072 11.532 ;
    END
  END w0_wd_in[1]
  PIN w0_wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 7.764 10.203 7.788 ;
    END
  END w0_wd_in[2]
  PIN w0_wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 11.508 10.203 11.532 ;
    END
  END w0_wd_in[3]
  PIN w0_wd_in[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 0.207 0.000 0.225 0.054 ;
    END
  END w0_wd_in[4]
  PIN w0_wd_in[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 1.395 0.000 1.413 0.054 ;
    END
  END w0_wd_in[5]
  PIN w0_wd_in[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.583 0.000 2.601 0.054 ;
    END
  END w0_wd_in[6]
  PIN r0_rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.771 0.000 3.789 0.054 ;
    END
  END r0_rd_out[0]
  PIN r0_rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.959 0.000 4.977 0.054 ;
    END
  END r0_rd_out[1]
  PIN r0_rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.147 0.000 6.165 0.054 ;
    END
  END r0_rd_out[2]
  PIN r0_rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.335 0.000 7.353 0.054 ;
    END
  END r0_rd_out[3]
  PIN r0_rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 2.367 45.909 2.385 45.963 ;
    END
  END r0_rd_out[4]
  PIN r0_rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.087 45.909 3.105 45.963 ;
    END
  END r0_rd_out[5]
  PIN r0_rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 3.807 45.909 3.825 45.963 ;
    END
  END r0_rd_out[6]
  PIN w0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.252 0.072 15.276 ;
    END
  END w0_addr_in[0]
  PIN w0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.996 0.072 19.020 ;
    END
  END w0_addr_in[1]
  PIN w0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.740 0.072 22.764 ;
    END
  END w0_addr_in[2]
  PIN w0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.484 0.072 26.508 ;
    END
  END w0_addr_in[3]
  PIN w0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 15.252 10.203 15.276 ;
    END
  END w0_addr_in[4]
  PIN w0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 18.996 10.203 19.020 ;
    END
  END w0_addr_in[5]
  PIN w0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 22.740 10.203 22.764 ;
    END
  END w0_addr_in[6]
  PIN w0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 26.484 10.203 26.508 ;
    END
  END w0_addr_in[7]
  PIN r0_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.228 0.072 30.252 ;
    END
  END r0_addr_in[0]
  PIN r0_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.972 0.072 33.996 ;
    END
  END r0_addr_in[1]
  PIN r0_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.716 0.072 37.740 ;
    END
  END r0_addr_in[2]
  PIN r0_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.460 0.072 41.484 ;
    END
  END r0_addr_in[3]
  PIN r0_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 30.228 10.203 30.252 ;
    END
  END r0_addr_in[4]
  PIN r0_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 33.972 10.203 33.996 ;
    END
  END r0_addr_in[5]
  PIN r0_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 37.716 10.203 37.740 ;
    END
  END r0_addr_in[6]
  PIN r0_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 10.131 41.460 10.203 41.484 ;
    END
  END r0_addr_in[7]
  PIN w0_we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.527 45.909 4.545 45.963 ;
    END
  END w0_we_in
  PIN w0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.247 45.909 5.265 45.963 ;
    END
  END w0_ce_in
  PIN w0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 5.967 45.909 5.985 45.963 ;
    END
  END w0_clk
  PIN r0_ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.687 45.909 6.705 45.963 ;
    END
  END r0_ce_in
  PIN r0_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 7.407 45.909 7.425 45.963 ;
    END
  END r0_clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
      RECT 0.216 13.296 9.987 13.392 ;
      RECT 0.216 14.064 9.987 14.160 ;
      RECT 0.216 14.832 9.987 14.928 ;
      RECT 0.216 15.600 9.987 15.696 ;
      RECT 0.216 16.368 9.987 16.464 ;
      RECT 0.216 17.136 9.987 17.232 ;
      RECT 0.216 17.904 9.987 18.000 ;
      RECT 0.216 18.672 9.987 18.768 ;
      RECT 0.216 19.440 9.987 19.536 ;
      RECT 0.216 20.208 9.987 20.304 ;
      RECT 0.216 20.976 9.987 21.072 ;
      RECT 0.216 21.744 9.987 21.840 ;
      RECT 0.216 22.512 9.987 22.608 ;
      RECT 0.216 23.280 9.987 23.376 ;
      RECT 0.216 24.048 9.987 24.144 ;
      RECT 0.216 24.816 9.987 24.912 ;
      RECT 0.216 25.584 9.987 25.680 ;
      RECT 0.216 26.352 9.987 26.448 ;
      RECT 0.216 27.120 9.987 27.216 ;
      RECT 0.216 27.888 9.987 27.984 ;
      RECT 0.216 28.656 9.987 28.752 ;
      RECT 0.216 29.424 9.987 29.520 ;
      RECT 0.216 30.192 9.987 30.288 ;
      RECT 0.216 30.960 9.987 31.056 ;
      RECT 0.216 31.728 9.987 31.824 ;
      RECT 0.216 32.496 9.987 32.592 ;
      RECT 0.216 33.264 9.987 33.360 ;
      RECT 0.216 34.032 9.987 34.128 ;
      RECT 0.216 34.800 9.987 34.896 ;
      RECT 0.216 35.568 9.987 35.664 ;
      RECT 0.216 36.336 9.987 36.432 ;
      RECT 0.216 37.104 9.987 37.200 ;
      RECT 0.216 37.872 9.987 37.968 ;
      RECT 0.216 38.640 9.987 38.736 ;
      RECT 0.216 39.408 9.987 39.504 ;
      RECT 0.216 40.176 9.987 40.272 ;
      RECT 0.216 40.944 9.987 41.040 ;
      RECT 0.216 41.712 9.987 41.808 ;
      RECT 0.216 42.480 9.987 42.576 ;
      RECT 0.216 43.248 9.987 43.344 ;
      RECT 0.216 44.016 9.987 44.112 ;
      RECT 0.216 44.784 9.987 44.880 ;
      RECT 0.216 45.552 9.987 45.648 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.216 0.240 9.987 0.336 ;
      RECT 0.216 1.008 9.987 1.104 ;
      RECT 0.216 1.776 9.987 1.872 ;
      RECT 0.216 2.544 9.987 2.640 ;
      RECT 0.216 3.312 9.987 3.408 ;
      RECT 0.216 4.080 9.987 4.176 ;
      RECT 0.216 4.848 9.987 4.944 ;
      RECT 0.216 5.616 9.987 5.712 ;
      RECT 0.216 6.384 9.987 6.480 ;
      RECT 0.216 7.152 9.987 7.248 ;
      RECT 0.216 7.920 9.987 8.016 ;
      RECT 0.216 8.688 9.987 8.784 ;
      RECT 0.216 9.456 9.987 9.552 ;
      RECT 0.216 10.224 9.987 10.320 ;
      RECT 0.216 10.992 9.987 11.088 ;
      RECT 0.216 11.760 9.987 11.856 ;
      RECT 0.216 12.528 9.987 12.624 ;
      RECT 0.216 13.296 9.987 13.392 ;
      RECT 0.216 14.064 9.987 14.160 ;
      RECT 0.216 14.832 9.987 14.928 ;
      RECT 0.216 15.600 9.987 15.696 ;
      RECT 0.216 16.368 9.987 16.464 ;
      RECT 0.216 17.136 9.987 17.232 ;
      RECT 0.216 17.904 9.987 18.000 ;
      RECT 0.216 18.672 9.987 18.768 ;
      RECT 0.216 19.440 9.987 19.536 ;
      RECT 0.216 20.208 9.987 20.304 ;
      RECT 0.216 20.976 9.987 21.072 ;
      RECT 0.216 21.744 9.987 21.840 ;
      RECT 0.216 22.512 9.987 22.608 ;
      RECT 0.216 23.280 9.987 23.376 ;
      RECT 0.216 24.048 9.987 24.144 ;
      RECT 0.216 24.816 9.987 24.912 ;
      RECT 0.216 25.584 9.987 25.680 ;
      RECT 0.216 26.352 9.987 26.448 ;
      RECT 0.216 27.120 9.987 27.216 ;
      RECT 0.216 27.888 9.987 27.984 ;
      RECT 0.216 28.656 9.987 28.752 ;
      RECT 0.216 29.424 9.987 29.520 ;
      RECT 0.216 30.192 9.987 30.288 ;
      RECT 0.216 30.960 9.987 31.056 ;
      RECT 0.216 31.728 9.987 31.824 ;
      RECT 0.216 32.496 9.987 32.592 ;
      RECT 0.216 33.264 9.987 33.360 ;
      RECT 0.216 34.032 9.987 34.128 ;
      RECT 0.216 34.800 9.987 34.896 ;
      RECT 0.216 35.568 9.987 35.664 ;
      RECT 0.216 36.336 9.987 36.432 ;
      RECT 0.216 37.104 9.987 37.200 ;
      RECT 0.216 37.872 9.987 37.968 ;
      RECT 0.216 38.640 9.987 38.736 ;
      RECT 0.216 39.408 9.987 39.504 ;
      RECT 0.216 40.176 9.987 40.272 ;
      RECT 0.216 40.944 9.987 41.040 ;
      RECT 0.216 41.712 9.987 41.808 ;
      RECT 0.216 42.480 9.987 42.576 ;
      RECT 0.216 43.248 9.987 43.344 ;
      RECT 0.216 44.016 9.987 44.112 ;
      RECT 0.216 44.784 9.987 44.880 ;
      RECT 0.216 45.552 9.987 45.648 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 10.203 45.963 ;
    LAYER M2 ;
    RECT 0 0 10.203 45.963 ;
    LAYER M3 ;
    RECT 0 0 10.203 45.963 ;
    LAYER M4 ;
    RECT 0 0 10.203 45.963 ;
  END
END fakeram_7x256_1r1w

END LIBRARY
